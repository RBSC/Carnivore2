-- megafunction wizard: %LPM_RAM_DQ%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_ram_dq 

-- ============================================================
-- File Name: ram.vhd
-- Megafunction Name(s):
--                      lpm_ram_dq
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--      Copyright (C) 1988-2000 Altera Corporation

--      Any megafunction design, and related net list (encrypted or decrypted),
--      support information, device programming or simulation file, and any other
--      associated documentation or information provided by Altera or a partner
--      under Altera's Megafunction Partnership Program may be used only to
--      program PLD devices (but not masked PLD devices) from Altera.  Any other
--      use of such megafunction design, net list, support information, device
--      programming or simulation file, or any other related documentation or
--      information is prohibited for any other purpose, including, but not
--      limited to modification, reverse engineering, de-compiling, or use with
--      any other silicon devices, unless such use is explicitly licensed under
--      a separate agreement with Altera or a megafunction partner.  Title to
--      the intellectual property, including patents, copyrights, trademarks,
--      trade secrets, or maskworks, embodied in any such megafunction design,
--      net list, support information, device programming or simulation file, or
--      any other related documentation or information provided by Altera or a
--      megafunction partner, remains with Altera, the megafunction partner, or
--      their respective licensors.  No other licenses, including any licenses
--      needed under any third party's intellectual property, are provided herein.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY ram IS
        PORT
        (
                address         : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                inclock         : IN STD_LOGIC ;
                we              : IN STD_LOGIC  := '1';
                data            : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                q               : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );
END ram;


ARCHITECTURE SYN OF ram IS

        SIGNAL sub_wire0        : STD_LOGIC_VECTOR (7 DOWNTO 0);



        COMPONENT lpm_ram_dq
        GENERIC (
                LPM_WIDTH               : NATURAL;
                LPM_WIDTHAD             : NATURAL;
                LPM_INDATA              : STRING;
                LPM_ADDRESS_CONTROL             : STRING;
                LPM_OUTDATA             : STRING;
                LPM_HINT                : STRING
        );
        PORT (
                        address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                        inclock : IN STD_LOGIC ;
                        q       : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                        data    : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                        we      : IN STD_LOGIC 
        );
        END COMPONENT;

BEGIN
        q    <= sub_wire0(7 DOWNTO 0);

        lpm_ram_dq_component : lpm_ram_dq
        GENERIC MAP (
                LPM_WIDTH => 8,
                LPM_WIDTHAD => 8,
                LPM_INDATA => "REGISTERED",
                LPM_ADDRESS_CONTROL => "REGISTERED",
                LPM_OUTDATA => "UNREGISTERED",
                LPM_HINT => "USE_EAB"
        )
        PORT MAP (
                address => address,
                inclock => inclock,
                data => data,
                we => we,
                q => sub_wire0
        );



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: WidthData NUMERIC "8"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "8"
-- Retrieval info: PRIVATE: RegData NUMERIC "1"
-- Retrieval info: PRIVATE: RegAdd NUMERIC "1"
-- Retrieval info: PRIVATE: OutputRegistered NUMERIC "0"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: UseLCs NUMERIC "0"
-- Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_WIDTHAD NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_INDATA STRING "REGISTERED"
-- Retrieval info: CONSTANT: LPM_ADDRESS_CONTROL STRING "REGISTERED"
-- Retrieval info: CONSTANT: LPM_OUTDATA STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "USE_EAB=ON"
-- Retrieval info: USED_PORT: address 0 0 8 0 INPUT NODEFVAL address[7..0]
-- Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT NODEFVAL inclock
-- Retrieval info: USED_PORT: we 0 0 0 0 INPUT VCC we
-- Retrieval info: USED_PORT: q 0 0 8 0 OUTPUT NODEFVAL q[7..0]
-- Retrieval info: USED_PORT: data 0 0 8 0 INPUT NODEFVAL data[7..0]
-- Retrieval info: CONNECT: @address 0 0 8 0 address 0 0 8 0
-- Retrieval info: CONNECT: @inclock 0 0 0 0 inclock 0 0 0 0
-- Retrieval info: CONNECT: @we 0 0 0 0 we 0 0 0 0
-- Retrieval info: CONNECT: q 0 0 8 0 @q 0 0 8 0
-- Retrieval info: CONNECT: @data 0 0 8 0 data 0 0 8 0
